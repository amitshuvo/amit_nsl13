class main
    bit a;
    bit b;
endclass: main
